INT_OSC_inst : INT_OSC PORT MAP (
		oscena	 => oscena_sig,
		osc	 => osc_sig
	);
