-- i2c_CORE.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity i2c_CORE is
	port (
		a0           : in    std_logic := '0'; --           a0.a0
		a1           : in    std_logic := '0'; --           a1.a1
		a2           : in    std_logic := '0'; --           a2.a2
		global_reset : in    std_logic := '0'; -- global_reset.global_reset
		osc          : out   std_logic;        --          osc.osc
		scl          : inout std_logic := '0'; --          scl.scl
		sda          : inout std_logic := '0'  --          sda.sda
	);
end entity i2c_CORE;

architecture rtl of i2c_CORE is
	component i2c_CORE_ufm_i2c_0 is
		port (
			a0           : in    std_logic := 'X'; -- a0
			a1           : in    std_logic := 'X'; -- a1
			a2           : in    std_logic := 'X'; -- a2
			scl          : inout std_logic := 'X'; -- scl
			sda          : inout std_logic := 'X'; -- sda
			global_reset : in    std_logic := 'X'; -- global_reset
			osc          : out   std_logic         -- osc
		);
	end component i2c_CORE_ufm_i2c_0;

begin

	ufm_i2c_0 : component i2c_CORE_ufm_i2c_0
		port map (
			a0           => a0,           --           a0.a0
			a1           => a1,           --           a1.a1
			a2           => a2,           --           a2.a2
			scl          => scl,          --          scl.scl
			sda          => sda,          --          sda.sda
			global_reset => global_reset, -- global_reset.global_reset
			osc          => osc           --          osc.osc
		);

end architecture rtl; -- of i2c_CORE
